module imem(input logic [31:0] a,
output logic [31:0] rd);
logic [31:0] RAM[255:0];// cambiar para progrs largos
initial
$readmemh("riscvtest.txt",RAM);
assign rd = RAM[a[31:2]]; // word aligned
endmodule
//AltGr +   ~

module dmem(input logic clk, we,input logic [31:0] a,
wd,output logic [31:0] rd,
input logic cs);

logic [31:0] RAM[255:0];//data=32bits dir=0-63(64localidades de 32 bits)
logic [31:0]ax;
assign ax=a & 32'H0FFFFFFF;
assign rd =cs? 32'bz : RAM[ax[31:2]]; // word aligned

always_ff @(posedge clk)
if(!cs)begin // habilita con oe=0
    if (we)RAM[ax[31:2]] <= wd; 
        end

initial begin
/*
        RAM[0] =~ 32'hC6C6C600;//fila 13,9,5,1
        RAM[1] =~ 32'hFEC6C6FE;//fila 14,10,6,2
        RAM[2] =~ 32'hFEC6C6FE;//fila 15,11,7,3
        RAM[3] =~ 32'h00C6C6C6;//fila 16,12,8,4

        RAM[4] =~ 32'h10011001;//fila 13,9,5,1 BLOCK8_0
        RAM[5] =~ 32'h20022002;//fila 14,10,6,2 BLOCK8_0
        RAM[6] =~ 32'h40044004;//fila 15,11,7,3 BLOCK8_0
        RAM[7] =~ 32'h80088008;//fila 16,12,8,4 BLOCK8_0

         RAM[8] =~ 32'h1c1c1c3c;//fila 13,9,5,1 BLOCK8_0
         RAM[9] =~ 32'h7f1c1c3c;//fila 14,10,6,2 BLOCK8_0
        RAM[10] =~ 32'h7f1c1c3c;//fila 15,11,7,3 BLOCK8_0
        RAM[11] =~ 32'h7f1c1c1c;//fila 16,12,8,4 BLOCK8_0

        RAM[12] =~ 32'h707F077F;//fila 13,9,5,1 BLOCK8_0
        RAM[13] =~ 32'h7F7F077F;//fila 14,10,6,2 BLOCK8_0
        RAM[14] =~ 32'h7F70077F;//fila 15,11,7,3 BLOCK8_0
        RAM[15] =~ 32'h7F707F07;//fila 16,12,8,4 BLOCK8_0
*/
RAM[0] = ~32'h00020000;
RAM[1] = ~32'h00000000;
RAM[2] = ~32'h00000000;
RAM[3] = ~32'h00000100;
RAM[4] = ~32'h243C7E00;
RAM[5] = ~32'h423C7E42;
RAM[6] = ~32'h423C7E7E;
RAM[7] = ~32'h0024BD5A;
RAM[8] = ~32'h00400000;
RAM[9] = ~32'h00000000;
RAM[10] = ~32'h00000000;
RAM[11] = ~32'h00008000;
RAM[12] = ~32'h00000000;
RAM[13] = ~32'h00000000;
RAM[14] = ~32'h00000000;
RAM[15] = ~32'h00000000;
RAM[16] = ~32'h00010000;
RAM[17] = ~32'h00000000;
RAM[18] = ~32'h00000000;
RAM[19] = ~32'h00000000;
RAM[20] = ~32'h121E3F00;
RAM[21] = ~32'h121E3F21;
RAM[22] = ~32'h121E3F3F;
RAM[23] = ~32'h0012DE2D;
RAM[24] = ~32'h00200000;
RAM[25] = ~32'h00000000;
RAM[26] = ~32'h00000000;
RAM[27] = ~32'h0000C000;
RAM[28] = ~32'h00000000;
RAM[29] = ~32'h00000000;
RAM[30] = ~32'h00000000;
RAM[31] = ~32'h00000000;
RAM[32] = ~32'h00000000;
RAM[33] = ~32'h00000000;
RAM[34] = ~32'h00000000;
RAM[35] = ~32'h00000000;
RAM[36] = ~32'h091F1F00;
RAM[37] = ~32'h100F1F10;
RAM[38] = ~32'h100F1F1F;
RAM[39] = ~32'h00091F16;
RAM[40] = ~32'h00808000;
RAM[41] = ~32'h80008080;
RAM[42] = ~32'h80008080;
RAM[43] = ~32'h00008080;
RAM[44] = ~32'h00000000;
RAM[45] = ~32'h00000000;
RAM[46] = ~32'h00000000;
RAM[47] = ~32'h00000000;
RAM[48] = ~32'h00000000;
RAM[49] = ~32'h00000000;
RAM[50] = ~32'h00000000;
RAM[51] = ~32'h00000000;
RAM[52] = ~32'h040F0F00;
RAM[53] = ~32'h04070F08;
RAM[54] = ~32'h04070F0F;
RAM[55] = ~32'h00040F0B;
RAM[56] = ~32'h80C0C000;
RAM[57] = ~32'h8080C040;
RAM[58] = ~32'h8080C0C0;
RAM[59] = ~32'h0080C040;
RAM[60] = ~32'h00000000;
RAM[61] = ~32'h00000000;
RAM[62] = ~32'h00000000;
RAM[63] = ~32'h00000000;
RAM[64] = ~32'h00000000;
RAM[65] = ~32'h00000000;
RAM[66] = ~32'h00000000;
RAM[67] = ~32'h00000000;
RAM[68] = ~32'h02230700;
RAM[69] = ~32'h04030704;
RAM[70] = ~32'h04030707;
RAM[71] = ~32'h00021B05;
RAM[72] = ~32'h40C4E000;
RAM[73] = ~32'h20C0E020;
RAM[74] = ~32'h20C0E0E0;
RAM[75] = ~32'h0040D8A0;
RAM[76] = ~32'h00000000;
RAM[77] = ~32'h00000000;
RAM[78] = ~32'h00000000;
RAM[79] = ~32'h00000000;
RAM[80] = ~32'h00000000;
RAM[81] = ~32'h00000000;
RAM[82] = ~32'h00000000;
RAM[83] = ~32'h00000000;
RAM[84] = ~32'h01110300;
RAM[85] = ~32'h01010302;
RAM[86] = ~32'h01010303;
RAM[87] = ~32'h00010D02;
RAM[88] = ~32'h20E2F000;
RAM[89] = ~32'h20E0F010;
RAM[90] = ~32'h20E0F0F0;
RAM[91] = ~32'h0020ECD0;
RAM[92] = ~32'h00000000;
RAM[93] = ~32'h00000000;
RAM[94] = ~32'h00000000;
RAM[95] = ~32'h00000000;
RAM[96] = ~32'h00000000;
RAM[97] = ~32'h00000000;
RAM[98] = ~32'h00000000;
RAM[99] = ~32'h00000000;
RAM[100] = ~32'h00010100;
RAM[101] = ~32'h01000101;
RAM[102] = ~32'h01000101;
RAM[103] = ~32'h00000101;
RAM[104] = ~32'h90F8F800;
RAM[105] = ~32'h08F0F808;
RAM[106] = ~32'h08F0F8F8;
RAM[107] = ~32'h0090F868;
RAM[108] = ~32'h00000000;
RAM[109] = ~32'h00000000;
RAM[110] = ~32'h00000000;
RAM[111] = ~32'h00000000;
RAM[112] = ~32'h00000000;
RAM[113] = ~32'h00000000;
RAM[114] = ~32'h00000000;
RAM[115] = ~32'h00000000;
RAM[116] = ~32'h00000000;
RAM[117] = ~32'h00000000;
RAM[118] = ~32'h00000000;
RAM[119] = ~32'h00000000;
RAM[120] = ~32'h48FCFC00;
RAM[121] = ~32'h4878FC84;
RAM[122] = ~32'h4878FCFC;
RAM[123] = ~32'h0048FCB4;
RAM[124] = ~32'h00000000;
RAM[125] = ~32'h00000000;
RAM[126] = ~32'h00000000;
RAM[127] = ~32'h00000000;
RAM[128] = ~32'h00000000;
RAM[129] = ~32'h00000000;
RAM[130] = ~32'h00000000;
RAM[131] = ~32'h00000000;
RAM[132] = ~32'h00020000;
RAM[133] = ~32'h00000000;
RAM[134] = ~32'h00000000;
RAM[135] = ~32'h00000100;
RAM[136] = ~32'h243C7E00;
RAM[137] = ~32'h423C7E42;
RAM[138] = ~32'h423C7E7E;
RAM[139] = ~32'h0024BD5A;
RAM[140] = ~32'h00400000;
RAM[141] = ~32'h00000000;
RAM[142] = ~32'h00000000;
RAM[143] = ~32'h00008000;
RAM[144] = ~32'h00000000;
RAM[145] = ~32'h00000000;
RAM[146] = ~32'h00000000;
RAM[147] = ~32'h00000000;
RAM[148] = ~32'h00010000;
RAM[149] = ~32'h00000000;
RAM[150] = ~32'h00000000;
RAM[151] = ~32'h00000000;
RAM[152] = ~32'h121E3F00;
RAM[153] = ~32'h121E3F21;
RAM[154] = ~32'h121E3F3F;
RAM[155] = ~32'h0012DE2D;
RAM[156] = ~32'h00200000;
RAM[157] = ~32'h00000000;
RAM[158] = ~32'h00000000;
RAM[159] = ~32'h0000C000;
RAM[160] = ~32'h00000000;
RAM[161] = ~32'h00000000;
RAM[162] = ~32'h00000000;
RAM[163] = ~32'h00000000;
RAM[164] = ~32'h00000000;
RAM[165] = ~32'h00000000;
RAM[166] = ~32'h00000000;
RAM[167] = ~32'h00000000;
RAM[168] = ~32'h091F1F00;
RAM[169] = ~32'h100F1F10;
RAM[170] = ~32'h100F1F1F;
RAM[171] = ~32'h00091F16;
RAM[172] = ~32'h00808000;
RAM[173] = ~32'h80008080;
RAM[174] = ~32'h80008080;
RAM[175] = ~32'h00008080;
RAM[176] = ~32'h00000000;
RAM[177] = ~32'h00000000;
RAM[178] = ~32'h00000000;
RAM[179] = ~32'h00000000;
RAM[180] = ~32'h00000000;
RAM[181] = ~32'h00000000;
RAM[182] = ~32'h00000000;
RAM[183] = ~32'h00000000;
RAM[184] = ~32'h040F0F00;
RAM[185] = ~32'h04070F08;
RAM[186] = ~32'h04070F0F;
RAM[187] = ~32'h00040F0B;
RAM[188] = ~32'h80C0C000;
RAM[189] = ~32'h8080C040;
RAM[190] = ~32'h8080C0C0;
RAM[191] = ~32'h0080C040;
RAM[192] = ~32'h00000000;
RAM[193] = ~32'h00000000;
RAM[194] = ~32'h00000000;
RAM[195] = ~32'h00000000;
RAM[196] = ~32'h00000000;
RAM[197] = ~32'h00000000;
RAM[198] = ~32'h00000000;
RAM[199] = ~32'h00000000;
RAM[200] = ~32'h02230700;
RAM[201] = ~32'h04030704;
RAM[202] = ~32'h04030707;
RAM[203] = ~32'h00021B05;
RAM[204] = ~32'h40C4E000;
RAM[205] = ~32'h20C0E020;
RAM[206] = ~32'h20C0E0E0;
RAM[207] = ~32'h0040D8A0;
RAM[208] = ~32'h00000000;
RAM[209] = ~32'h00000000;
RAM[210] = ~32'h00000000;
RAM[211] = ~32'h00000000;
RAM[212] = ~32'h00000000;
RAM[213] = ~32'h00000000;
RAM[214] = ~32'h00000000;
RAM[215] = ~32'h00000000;
RAM[216] = ~32'h01110300;
RAM[217] = ~32'h01010302;
RAM[218] = ~32'h01010303;
RAM[219] = ~32'h00010D02;
RAM[220] = ~32'h20E2F000;
RAM[221] = ~32'h20E0F010;
RAM[222] = ~32'h20E0F0F0;
RAM[223] = ~32'h0020ECD0;
RAM[224] = ~32'h00000000;
RAM[225] = ~32'h00000000;
RAM[226] = ~32'h00000000;
RAM[227] = ~32'h00000000;
RAM[228] = ~32'h00000000;
RAM[229] = ~32'h00000000;
RAM[230] = ~32'h00000000;
RAM[231] = ~32'h00000000;
RAM[232] = ~32'h00010100;
RAM[233] = ~32'h01000101;
RAM[234] = ~32'h01000101;
RAM[235] = ~32'h00000101;
RAM[236] = ~32'h90F8F800;
RAM[237] = ~32'h08F0F808;
RAM[238] = ~32'h08F0F8F8;
RAM[239] = ~32'h0090F868;
RAM[240] = ~32'h00000000;
RAM[241] = ~32'h00000000;
RAM[242] = ~32'h00000000;
RAM[243] = ~32'h00000000;
RAM[244] = ~32'h00000000;
RAM[245] = ~32'h00000000;
RAM[246] = ~32'h00000000;
RAM[247] = ~32'h00000000;
RAM[248] = ~32'h00000000;
RAM[249] = ~32'h00000000;
RAM[250] = ~32'h00000000;
RAM[251] = ~32'h00000000;
RAM[252] = ~32'h48FCFC00;
RAM[253] = ~32'h4878FC84;
RAM[254] = ~32'h4878FCFC;
RAM[255] = ~32'h0048FCB4;      // puedes continuar hasta mem[31]

end

endmodule


module rom_32X16_uu(input logic [7:0]dir, output logic [15:0]data);
logic [31:0]dir_uu[0:255];//[0:87]
initial begin // módulos para poner letras
//cer0
dir_uu[00]=32'H00000000;
dir_uu[01]=32'H00000000;
dir_uu[02]=32'H00000000;
dir_uu[03]=32'H00000000;

end
endmodule